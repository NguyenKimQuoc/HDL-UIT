library verilog;
use verilog.vl_types.all;
entity TestFmulti is
end TestFmulti;
