library verilog;
use verilog.vl_types.all;
entity TestModule is
end TestModule;
