library verilog;
use verilog.vl_types.all;
entity Counter_NBIT_vlg_vec_tst is
end Counter_NBIT_vlg_vec_tst;
