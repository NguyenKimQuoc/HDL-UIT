module queue(io, empty, full, reset_n, en, rw, clk);
  parameter N = 11;
  parameter M = 8;
  inout [7:0] io;
  
  input reset_n, en, rw, clk;
  output empty, full;
  wire [10:0] out_cnt1;
  wire [10:0] out_cnt2;
  wire [9:0] out_mux;
  wire rw_n, mux_ctrl, en_cnt1, en_cnt2, RWS, out_comparator;
  
  not n1(rw_n, rw);
  and a1(en_cnt1, en, rw_n);
  and a2(en_cnt2, en, rw);
  Counter cnt1(out_cnt1[10:0], 0, en_cnt1, reset_n, clk); //cnt 11  bit
  Counter cnt2(out_cnt2[10:0], 0, en_cnt2, reset_n, clk); 
  
  and a3(mux_ctrl, en, rw_n);
  Mux_2to1_10bit mux(out_mux[9:0], out_cnt2[9:0], out_cnt1[9:0], mux_ctrl);
  Comparator cmp(out_comparator, out_cnt2[9:0], out_cnt1[9:0]);
  and a4(RWS, en, rw);  
  
  RAM r(io, out_mux[9:0], RWS, en, 1);
  xor xx1(x1, out_cnt2[10], out_cnt1[10]);
  not n2(x1_n, x1);
  and a5(empty, x1_n, out_comparator);
  and a6(full, x1, out_comparator);
endmodule