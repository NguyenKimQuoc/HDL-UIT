library verilog;
use verilog.vl_types.all;
entity TestFdivider is
end TestFdivider;
