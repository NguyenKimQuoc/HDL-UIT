library verilog;
use verilog.vl_types.all;
entity Stack_vlg_vec_tst is
end Stack_vlg_vec_tst;
