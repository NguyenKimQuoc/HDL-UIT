library verilog;
use verilog.vl_types.all;
entity SRwPLtest is
end SRwPLtest;
