library verilog;
use verilog.vl_types.all;
entity tb_DFF is
end tb_DFF;
