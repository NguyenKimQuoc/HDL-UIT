library verilog;
use verilog.vl_types.all;
entity TestDegtoRad is
end TestDegtoRad;
