library verilog;
use verilog.vl_types.all;
entity tb_Counter_8BIT is
end tb_Counter_8BIT;
