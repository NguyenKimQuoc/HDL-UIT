library verilog;
use verilog.vl_types.all;
entity TestDecoder is
end TestDecoder;
